LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY part2 IS
PORT(SW :IN STD_LOGIC_VECTOR(17 DOWNTO 0);
	  LEDG :OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END part2;

ARCHITECTURE Behavior OF part2 IS
BEGIN
LEDG(7) <= (NOT SW(17) AND SW(16)) OR (SW(17) AND SW(15));
LEDG(6) <= (NOT SW(17) AND SW(14)) OR (SW(17) AND SW(13));
LEDG(5) <= (NOT SW(17) AND SW(12)) OR (SW(17) AND SW(11));
LEDG(4) <= (NOT SW(17) AND SW(10)) OR (SW(17) AND SW(9));
LEDG(3) <= (NOT SW(17) AND SW(8)) OR (SW(17) AND SW(7));
LEDG(2) <= (NOT SW(17) AND SW(6)) OR (SW(17) AND SW(5));
LEDG(1) <= (NOT SW(17) AND SW(4)) OR (SW(17) AND SW(3));
LEDG(0) <= (NOT SW(17) AND SW(2)) OR (SW(17) AND SW(1));
END Behavior;